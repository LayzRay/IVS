//Опишем дешифратор для вывода на индикаторы. За основу возьмём дешифратор из 2-ой лабораторной.

module DC (X, Y);

	input [3:0] X;
	output reg [6:0] Y;
	
	always @( X ) begin
	
		case( X[3:0] )	
		
				4'b0000:    Y <= 7'b1000_000; // 0
				4'b0001:	Y <= 7'b1111_001; // 1
				4'b0010:	Y <= 7'b0100_100; // 2
				4'b0011:	Y <= 7'b0110_000; // 3
				4'b0100:	Y <= 7'b0011_001; // 4
				4'b0101:	Y <= 7'b0010_010; // 5
				4'b0110:    Y <= 7'b0000_010; // 6
				4'b0111:	Y <= 7'b1111_000; // 7
				4'b1000:	Y <= 7'b0000_000; // 8
				4'b1001:	Y <= 7'b0010_000; // 9
				4'b1010:	Y <= 7'b0001_000; // A
				4'b1011:	Y <= 7'b0000_011; // B
				4'b1100:	Y <= 7'b1000_110; // C
				4'b1101:	Y <= 7'b0100_001; // D
				4'b1110:	Y <= 7'b0000_110; // E
				4'b1111:	Y <= 7'b0001_110; // F
					
				default:    Y <= 7'b1111_111;
				
			endcase
	
	end
	
endmodule


